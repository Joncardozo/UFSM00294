module BCD7Seg (
	input [3:0] num,
	output [7:0] code
);

	assign code = 
			 (num == 4'b0000) ? 8'b11000000 : // 0
			 (num == 4'b0001) ? 8'b11111001 : // 1
			 (num == 4'b0010) ? 8'b10100100 : // 2
			 (num == 4'b0011) ? 8'b10110000 : // 3 
			 (num == 4'b0100) ? 8'b10011001 : // 4
			 (num == 4'b0101) ? 8'b10010010 : // 5
			 (num == 4'b0110) ? 8'b10000010 : // 6
			 (num == 4'b0111) ? 8'b11111000 : // 7
			 (num == 4'b1000) ? 8'b10000000 : // 8
			 (num == 4'b1001) ? 8'b10010000 : // 9 
			 (num == 4'b1010) ? 8'b10001000 : // A
			 (num == 4'b1011) ? 8'b10000011 : // b
			 (num == 4'b1100) ? 8'b11000110 : // C
			 (num == 4'b1101) ? 8'b10100001 : // d
			 (num == 4'b1110) ? 8'b10000110 : // E
			 (num == 4'b1111) ? 8'b10001110 : // F
									 8'b11111111 ; // apagado (valor inválido)


endmodule